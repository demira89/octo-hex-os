conectix             ,�'�qemu  Wi2k     @H      @H  y   ���ݺ:o��N�7�%�N                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������conectix             ,�'�qemu  Wi2k     @H      @H  y   ���ݺ:o��N�7�%�N                                                                                                                                                                                                                                                                                                                                                                                                                                            